** Generated on: Nov  6 18:36:39 2022
** Design library name: work_VR
** Design cell name: zz_oa_telescopicNin
** Design view name: schematic

** Library name: work_VR
** Cell name: oa_telescopicNin
** View name: schematic

.subckt oa_telescopicNin ib25a ibb50a ibc200a vdda vin vip vo vssa

** Telescopic OpAmp

** Top devices
m3 net4 vbpw vdda vdda tsmc18dP L=180e-9 W=1.44e-6 AD=648e-15 AS=648e-15 PD=3.78e-6 PS=3.78e-6 M=16
m4 net5 vbpw vdda vdda tsmc18dP L=180e-9 W=1.44e-6 AD=648e-15 AS=648e-15 PD=3.78e-6 PS=3.78e-6 M=16

** L2 Cascode
m3c net7 vbpcw net4 vdda tsmc18dP L=180e-9 W=1.44e-6 AD=648e-15 AS=648e-15 PD=3.78e-6 PS=3.78e-6 M=16
m4c vo vbpcw net5 vdda tsmc18dP L=180e-9 W=1.44e-6 AD=648e-15 AS=648e-15 PD=3.78e-6 PS=3.78e-6 M=16

** L1 Cascode
m1c net7 ibc200a net3 vssa tsmc18dN L=180e-9 W=720e-9 AD=324e-15 AS=324e-15 PD=2.34e-6 PS=2.34e-6 M=5
m2c vo ibc200a net6 vssa tsmc18dN L=180e-9 W=720e-9 AD=324e-15 AS=324e-15 PD=2.34e-6 PS=2.34e-6 M=5

** Cascode FETs bias device
m1cb ibc200a ibc200a vt vssa tsmc18dN L=180e-9 W=720e-9 AD=324e-15 AS=324e-15 PD=2.34e-6 PS=2.34e-6 M=5

** Input FETs
m2 net6 vip vt vssa tsmc18dN L=180e-9 W=720e-9 AD=324e-15 AS=324e-15 PD=2.34e-6 PS=2.34e-6 M=5
m1 net3 vin vt vssa tsmc18dN L=180e-9 W=720e-9 AD=324e-15 AS=324e-15 PD=2.34e-6 PS=2.34e-6 M=5

** Tail and current miror devices
m5 vt ib25a vssa vssa tsmc18dN L=1.44e-6 W=5.58e-6 AD=2.511e-12 AS=2.511e-12 PD=12.06e-6 PS=12.06e-6 M=16
m6 ib25a ib25a vssa vssa tsmc18dN L=1.44e-6 W=5.58e-6 AD=2.511e-12 AS=2.511e-12 PD=12.06e-6 PS=12.06e-6 M=2


** Wide-swing current mirror

m3r net2 vbpcw vdda vdda tsmc18dP L=180e-9 W=1.44e-6 AD=648e-15 AS=648e-15 PD=3.78e-6 PS=3.78e-6 M=16
m3bw net1 vbpw vdda vdda tsmc18dP L=180e-9 W=1.44e-6 AD=648e-15 AS=648e-15 PD=3.78e-6 PS=3.78e-6 M=16
m3cbw vbpcw vbpcw net2 vdda tsmc18dP L=180e-9 W=1.44e-6 AD=648e-15 AS=648e-15 PD=3.78e-6 PS=3.78e-6 M=16
m3bwc vbpw vbpcw net1 vdda tsmc18dP L=180e-9 W=1.44e-6 AD=648e-15 AS=648e-15 PD=3.78e-6 PS=3.78e-6 M=16

.param l0 = 1.44e-6
.param w0 = 5.58e-6
.param m0 = 2

** Tail current devices L2
m8c vbpw ibb50a net12 vssa tsmc18dN L=1.44e-6 W=5.58e-6 AD=2.511e-12 AS=2.511e-12 PD=12.06e-6 PS=12.06e-6 M=2
m7c vbpcw ibb50a net10 vssa tsmc18dN L=1.44e-6 W=5.58e-6 AD=2.511e-12 AS=2.511e-12 PD=12.06e-6 PS=12.06e-6 M=2

** Tail current devices L1
m7 net10 vbn vssa vssa tsmc18dN L=1.44e-6 W=5.58e-6 AD=2.511e-12 AS=2.511e-12 PD=12.06e-6 PS=12.06e-6 M=2
m8 net12 vbn vssa vssa tsmc18dN L=1.44e-6 W=5.58e-6 AD=2.511e-12 AS=2.511e-12 PD=12.06e-6 PS=12.06e-6 M=2

** Current mirror leg
m0c ibb50a ibb50a vbn vssa tsmc18dN L=1.44e-6 W=5.58e-6 AD=2.511e-12 AS=2.511e-12 PD=12.06e-6 PS=12.06e-6 M=2
m0 vbn vbn vssa vssa tsmc18dN L=1.44e-6 W=5.58e-6 AD=2.511e-12 AS=2.511e-12 PD=12.06e-6 PS=12.06e-6 M=2

.ends oa_telescopicNin
** End of subcircuit definition.
